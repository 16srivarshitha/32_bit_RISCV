module Instruction_decode(

);
endmodule