module execute(
    
);
endmodule